module fbitcomparator(input [3:0] a,[3:0] b,output gt,lt,eq);
    assign gt = a[3]&(~b[3]) + (~(a[3]^b[3]))&a[2]&(~b[2]) + (~(a[3]^b[3]))&(~(a[2]^b[2]))&a[1]&(~b[1]) + (~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]^b[1]))&(a[0]&(~b[0]));

    assign lt= (~a[3])&b[3]+(~(a[3]^b[3]))&(~a[2]&b[2])+(~(a[3]^b[3]))&(~(a[2]^b[2]))&(~a[1])&b[1] + (~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]^b[1]))&((~a[0])&b[0]);

    assign eq = (~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]^b[1]))&(~(a[0]^b[0]));

endmodule


